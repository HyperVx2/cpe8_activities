CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 20 30 110 10
1140 84 1914 1007
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
1308 180 1421 277
76546066 256
0
6 Title:
5 Name:
0
0
0
32
13 Logic Switch~
5 252 54 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21872 270
2 5V
-6 -21 8 -13
2 V4
-6 -31 8 -23
1 D
-3 -31 4 -23
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
366 0 0
2
44973.9 1
0
13 Logic Switch~
5 171 54 0 1 11
0 22
0
0 0 21872 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
1 C
-3 -31 4 -23
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5762 0 0
2
44973.9 1
0
13 Logic Switch~
5 90 54 0 1 11
0 12
0
0 0 21872 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
1 B
-3 -32 4 -24
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4943 0 0
2
44973.9 0
0
13 Logic Switch~
5 54 54 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21872 270
2 5V
-6 -21 8 -13
2 V1
-6 -31 8 -23
1 A
-3 -32 4 -24
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3435 0 0
2
44973.9 0
0
9 CC 7-Seg~
183 639 108 0 18 19
10 9 10 8 7 6 5 4 26 27
1 1 1 1 0 1 1 2 2
0
0 0 21088 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 0 0 0 0
4 DISP
8705 0 0
2
44973.9 0
0
14 Logic Display~
6 576 675 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4331 0 0
2
44973.9 0
0
14 Logic Display~
6 576 621 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
787 0 0
2
44973.9 0
0
14 Logic Display~
6 576 549 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3655 0 0
2
44973.9 0
0
14 Logic Display~
6 576 486 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6682 0 0
2
44973.9 0
0
14 Logic Display~
6 576 396 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
582 0 0
2
44973.9 0
0
14 Logic Display~
6 576 306 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3125 0 0
2
44973.9 0
0
14 Logic Display~
6 576 153 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
5466 0 0
2
44973.9 0
0
8 4-In OR~
219 531 693 0 5 22
0 15 2 14 3 4
0
0 0 1136 0
4 4072
-14 -24 14 -16
3 U9A
-3 -25 18 -17
1 g
-2 -26 5 -18
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 9 0
1 U
52 0 0
2
44973.9 0
0
8 4-In OR~
219 531 639 0 5 22
0 17 16 2 3 5
0
0 0 1136 0
4 4072
-14 -24 14 -16
3 U8B
-3 -25 18 -17
1 f
-1 -27 6 -19
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 8 0
1 U
3898 0 0
2
44973.9 0
0
5 4081~
219 360 630 0 3 22
0 12 13 16
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U5D
-12 -25 9 -17
3 B~D
-13 -27 8 -19
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
9413 0 0
2
44973.9 0
0
5 4081~
219 360 684 0 3 22
0 12 11 2
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U5C
-12 -25 9 -17
3 B~C
-12 -25 9 -17
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
8576 0 0
2
44973.9 0
0
5 4071~
219 531 567 0 3 22
0 18 15 6
0
0 0 1136 0
4 4071
-7 -24 21 -16
3 U7B
-3 -25 18 -17
1 e
-1 -25 6 -17
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 7 0
1 U
622 0 0
2
44973.9 0
0
8 4-In OR~
219 531 504 0 5 22
0 20 18 15 19 7
0
0 0 1136 0
4 4072
-14 -24 14 -16
3 U8A
-3 -25 18 -17
1 d
-2 -27 5 -19
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 8 0
1 U
9152 0 0
2
44973.9 0
0
5 4071~
219 477 468 0 3 22
0 3 14 20
0
0 0 1136 0
4 4071
-7 -24 21 -16
3 U7A
-3 -25 18 -17
5 A+~BC
-4 -26 31 -18
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
783 0 0
2
44973.9 0
0
5 4073~
219 360 576 0 4 22
0 12 11 21 19
0
0 0 1136 0
4 4073
-7 -24 21 -16
3 U6A
-12 -25 9 -17
4 B~CD
-16 -26 12 -18
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 6 0
1 U
4262 0 0
2
44973.9 0
0
5 4081~
219 360 522 0 3 22
0 22 13 15
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U5B
-12 -25 9 -17
3 C~D
-11 -26 10 -18
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
6121 0 0
2
44973.9 0
0
5 4081~
219 360 468 0 3 22
0 23 22 14
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
3 ~BC
-12 -25 9 -17
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
3879 0 0
2
44973.9 0
0
8 3-In OR~
219 531 414 0 4 22
0 12 11 21 8
0
0 0 1136 0
4 4075
-14 -24 14 -16
3 U4A
-3 -25 18 -17
1 c
-3 -26 4 -18
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 4 0
1 U
7345 0 0
2
44973.9 0
0
8 4-In OR~
219 531 324 0 5 22
0 3 23 24 17 10
0
0 0 1136 0
4 4072
-14 -24 14 -16
3 U3B
-3 -25 18 -17
1 b
-2 -27 5 -19
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 3 0
1 U
3198 0 0
2
44973.9 0
0
5 4081~
219 360 378 0 3 22
0 11 13 17
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U2D
-12 -25 9 -17
4 ~C~D
-18 -26 10 -18
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
9849 0 0
2
44973.9 0
0
5 4081~
219 360 324 0 3 22
0 22 21 24
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U2C
-12 -25 9 -17
2 CD
-12 -26 2 -18
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
479 0 0
2
44973.9 0
0
8 4-In OR~
219 531 171 0 5 22
0 3 22 18 25 9
0
0 0 1136 0
4 4072
-14 -24 14 -16
3 U3A
-3 -25 18 -17
1 a
-3 -27 4 -19
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 3 0
1 U
3905 0 0
2
44973.9 0
0
5 4081~
219 360 243 0 3 22
0 12 21 25
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
2 BD
-9 -25 5 -17
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
4394 0 0
2
44973.9 0
0
5 4081~
219 360 180 0 3 22
0 23 13 18
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
4 ~B~D
-17 -25 11 -17
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
4391 0 0
2
44973.9 0
0
5 4049~
219 279 99 0 2 22
0 21 13
0
0 0 1136 270
4 4049
-7 -24 21 -16
3 U1C
16 -8 37 0
2 ~D
17 -8 31 0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 1 0
1 U
3681 0 0
2
44973.9 0
0
5 4049~
219 198 99 0 2 22
0 22 11
0
0 0 1136 270
4 4049
-7 -24 21 -16
3 U1B
16 -8 37 0
2 ~C
18 -8 32 0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 1 0
1 U
6466 0 0
2
44973.9 0
0
5 4049~
219 117 99 0 2 22
0 12 23
0
0 0 1136 270
4 4049
-7 -24 21 -16
3 U1A
16 -8 37 0
2 ~B
17 -8 31 0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
5230 0 0
2
44973.9 0
0
70
2 0 2 0 0 8192 0 13 0 0 26 3
514 689
471 689
471 644
1 0 3 0 0 12288 0 19 0 0 70 4
464 459
385 459
385 429
54 429
1 0 4 0 0 0 0 6 0 0 4 2
576 693
576 693
5 7 4 0 0 8320 0 13 5 0 0 3
564 693
654 693
654 144
1 0 5 0 0 0 0 7 0 0 6 2
576 639
576 639
5 6 5 0 0 8320 0 14 5 0 0 3
564 639
648 639
648 144
1 0 6 0 0 0 0 8 0 0 8 2
576 567
576 567
3 5 6 0 0 8320 0 17 5 0 0 3
564 567
642 567
642 144
1 0 7 0 0 0 0 9 0 0 10 2
576 504
576 504
5 4 7 0 0 8320 0 18 5 0 0 3
564 504
636 504
636 144
1 0 8 0 0 0 0 10 0 0 12 2
576 414
576 414
4 3 8 0 0 8320 0 23 5 0 0 3
564 414
630 414
630 144
1 0 9 0 0 4096 0 12 0 0 16 2
576 171
576 170
1 0 10 0 0 0 0 11 0 0 15 2
576 324
576 324
5 2 10 0 0 8320 0 24 5 0 0 3
564 324
624 324
624 144
5 1 9 0 0 8320 0 27 5 0 0 4
564 171
564 170
618 170
618 144
2 0 11 0 0 4096 0 16 0 0 62 2
336 693
201 693
1 0 12 0 0 4096 0 16 0 0 69 2
336 675
90 675
2 0 13 0 0 4096 0 15 0 0 21 2
336 639
282 639
1 0 12 0 0 0 0 15 0 0 69 2
336 621
90 621
2 0 13 0 0 4224 0 30 0 0 21 3
282 117
282 750
283 750
4 0 3 0 0 8192 0 13 0 0 70 3
514 707
514 724
54 724
0 3 14 0 0 4224 0 0 13 35 0 3
457 477
457 698
514 698
0 1 15 0 0 4224 0 0 13 32 0 3
451 509
451 680
514 680
4 0 3 0 0 0 0 14 0 0 70 4
514 653
399 653
399 708
54 708
3 3 2 0 0 4224 0 14 16 0 0 4
514 644
389 644
389 684
381 684
2 3 16 0 0 4224 0 14 15 0 0 4
514 635
389 635
389 630
381 630
1 0 17 0 0 8320 0 14 0 0 50 3
514 626
443 626
443 338
2 0 15 0 0 0 0 17 0 0 32 3
518 576
430 576
430 509
1 0 18 0 0 8320 0 17 0 0 57 3
518 558
421 558
421 176
4 4 19 0 0 4224 0 18 20 0 0 4
514 518
394 518
394 576
381 576
3 3 15 0 0 0 0 18 21 0 0 4
514 509
389 509
389 522
381 522
0 2 18 0 0 0 0 0 18 57 0 3
406 176
406 500
514 500
3 1 20 0 0 4224 0 19 18 0 0 3
510 468
510 491
514 491
2 3 14 0 0 0 0 19 22 0 0 4
464 477
389 477
389 468
381 468
3 0 21 0 0 4096 0 20 0 0 67 2
336 585
252 585
2 0 11 0 0 0 0 20 0 0 62 2
336 576
201 576
1 0 12 0 0 0 0 20 0 0 69 2
336 567
90 567
2 0 13 0 0 0 0 21 0 0 21 2
336 531
282 531
1 0 22 0 0 4096 0 21 0 0 68 2
336 513
171 513
2 0 22 0 0 0 0 22 0 0 68 2
336 477
171 477
1 0 23 0 0 4096 0 22 0 0 63 2
336 459
120 459
3 0 21 0 0 4096 0 23 0 0 67 4
518 423
257 423
257 424
252 424
2 0 11 0 0 4096 0 23 0 0 62 2
519 414
201 414
1 0 12 0 0 4096 0 23 0 0 69 2
518 405
90 405
2 0 13 0 0 0 0 25 0 0 21 2
336 387
282 387
1 0 11 0 0 0 0 25 0 0 62 2
336 369
201 369
2 0 21 0 0 0 0 26 0 0 67 4
336 333
257 333
257 334
252 334
1 0 22 0 0 0 0 26 0 0 68 2
336 315
171 315
4 3 17 0 0 0 0 24 25 0 0 4
514 338
389 338
389 378
381 378
3 3 24 0 0 4224 0 24 26 0 0 4
514 329
389 329
389 324
381 324
2 0 23 0 0 12288 0 24 0 0 63 4
514 320
505 320
505 290
120 290
1 0 3 0 0 0 0 24 0 0 70 4
514 311
512 311
512 276
54 276
2 0 21 0 0 0 0 28 0 0 67 2
336 252
252 252
1 0 12 0 0 0 0 28 0 0 69 2
336 234
90 234
4 3 25 0 0 8320 0 27 28 0 0 5
514 185
514 196
396 196
396 243
381 243
3 3 18 0 0 0 0 27 29 0 0 4
514 176
389 176
389 180
381 180
2 0 22 0 0 12288 0 27 0 0 68 4
514 167
505 167
505 149
171 149
1 0 3 0 0 0 0 27 0 0 70 3
514 158
514 141
54 141
2 0 13 0 0 0 0 29 0 0 21 4
336 189
287 189
287 190
282 190
1 0 23 0 0 0 0 29 0 0 63 2
336 171
120 171
2 0 11 0 0 4224 0 31 0 0 0 2
201 117
201 755
2 0 23 0 0 4224 0 32 0 0 0 2
120 117
120 757
1 0 21 0 0 0 0 30 0 0 67 3
282 81
282 77
252 77
1 0 12 0 0 0 0 32 0 0 69 3
120 81
120 77
90 77
1 0 22 0 0 0 0 31 0 0 68 3
201 81
201 77
171 77
1 0 21 0 0 4224 0 1 0 0 0 2
252 66
252 754
1 0 22 0 0 4224 0 2 0 0 0 2
171 66
171 755
1 0 12 0 0 4224 0 3 0 0 0 2
90 66
90 757
1 0 3 0 0 4224 0 4 0 0 0 2
54 66
54 758
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
