CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 1 2 1
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 256
0
6 Title:
5 Name:
0
0
0
10
13 Logic Switch~
5 180 63 0 1 11
0 10
0
0 0 21872 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
1 C
-3 -30 4 -22
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4747 0 0
2
44974.4 1
0
13 Logic Switch~
5 108 63 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21872 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
1 B
-3 -31 4 -23
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
972 0 0
2
44974.4 0
0
13 Logic Switch~
5 27 63 0 1 11
0 8
0
0 0 21872 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
1 A
-4 -31 3 -23
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3472 0 0
2
44974.4 0
0
14 Logic Display~
6 405 144 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9998 0 0
2
44974.4 0
0
5 4071~
219 351 162 0 3 22
0 4 3 2
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U3A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
3536 0 0
2
44974.4 0
0
5 4081~
219 279 189 0 3 22
0 6 5 3
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
4 ~A~C
-16 -26 12 -18
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
4597 0 0
2
44974.4 0
0
5 4081~
219 279 135 0 3 22
0 6 7 4
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U2A
-12 -25 9 -17
4 ~A~B
-17 -25 11 -17
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
3835 0 0
2
44974.4 0
0
5 4049~
219 55 99 0 2 22
0 8 6
0
0 0 1136 270
4 4049
-7 -24 21 -16
3 U1C
16 -8 37 0
2 ~A
16 -8 30 0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 1 0
1 U
3670 0 0
2
44974.4 0
0
5 4049~
219 207 99 0 2 22
0 10 5
0
0 0 1136 270
4 4049
-7 -24 21 -16
3 U1B
16 -8 37 0
2 ~C
17 -8 31 0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 1 0
1 U
5616 0 0
2
44974.4 0
0
5 4049~
219 135 99 0 2 22
0 9 7
0
0 0 1136 270
4 4049
-7 -24 21 -16
3 U1A
16 -8 37 0
2 ~B
16 -8 30 0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
9323 0 0
2
44974.4 0
0
13
3 1 2 0 0 4224 0 5 4 0 0 2
384 162
405 162
2 3 3 0 0 4224 0 5 6 0 0 4
338 171
308 171
308 189
300 189
1 3 4 0 0 4224 0 5 7 0 0 4
338 153
308 153
308 135
300 135
2 0 5 0 0 4096 0 6 0 0 10 2
255 198
210 198
1 0 6 0 0 4224 0 6 0 0 8 2
255 180
58 180
2 0 7 0 0 4224 0 7 0 0 9 2
255 144
138 144
1 0 6 0 0 0 0 7 0 0 8 2
255 126
58 126
2 0 6 0 0 0 0 8 0 0 0 2
58 117
58 225
2 0 7 0 0 0 0 10 0 0 0 2
138 117
138 225
2 0 5 0 0 4224 0 9 0 0 0 2
210 117
210 225
1 1 8 0 0 8320 0 8 3 0 0 4
58 81
58 80
27 80
27 75
1 1 9 0 0 8320 0 10 2 0 0 4
138 81
138 80
108 80
108 75
1 1 10 0 0 8336 0 9 1 0 0 4
210 81
210 80
180 80
180 75
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
