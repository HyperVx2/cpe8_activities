CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
76546066 256
0
2 

2 

0
0
0
32
13 Logic Switch~
5 405 68 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21872 270
2 5V
-5 -33 9 -25
2 V4
-6 -26 8 -18
1 D
-3 -21 4 -13
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5636 0 0
2
44973.7 0
0
13 Logic Switch~
5 224 69 0 1 11
0 16
0
0 0 21872 270
2 0V
-6 -31 8 -23
2 V2
-6 -26 8 -18
1 B
-3 -21 4 -13
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
327 0 0
2
44973.7 1
0
13 Logic Switch~
5 308 68 0 1 11
0 22
0
0 0 21872 270
2 0V
-5 -33 9 -25
2 V3
-6 -26 8 -18
1 C
-3 -21 4 -13
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9233 0 0
2
44973.7 2
0
13 Logic Switch~
5 138 70 0 10 11
0 14 0 0 0 0 0 0 0 0
1
0
0 0 21872 270
2 5V
-6 -31 8 -23
2 V1
-6 -26 8 -18
1 A
-3 -18 4 -10
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3875 0 0
2
44973.7 3
0
5 4071~
219 664 655 0 3 22
0 4 6 5
0
0 0 1136 0
0
4 U10B
-6 -25 22 -17
12 4 terms+B~CD
-43 -31 41 -23
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 10 0
1 U
9991 0 0
2
44973.7 0
0
9 CC 7-Seg~
183 990 117 0 18 19
10 12 11 10 9 5 8 7 26 27
1 1 1 1 0 1 1 2 2
0
0 0 21088 0
6 BLUECC
13 -41 55 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3221 0 0
2
5.90066e-315 0
0
8 4-In OR~
219 665 756 0 5 22
0 14 2 19 18 8
0
0 0 1136 0
4 4072
-14 -24 14 -16
3 U4A
-3 -25 18 -17
1 f
-8 -29 -1 -21
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
8874 0 0
2
5.90066e-315 0
0
5 4071~
219 675 522 0 3 22
0 21 20 9
0
0 0 1136 0
0
4 U10A
-6 -25 22 -17
12 4 terms+B~CD
-43 -31 41 -23
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 10 0
1 U
7400 0 0
2
5.90066e-315 0
0
8 4-In OR~
219 675 414 0 5 22
0 14 16 17 3 10
0
0 0 1136 0
4 4072
-14 -24 14 -16
3 U9A
-3 -25 18 -17
1 c
-8 -29 -1 -21
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 9 0
1 U
3623 0 0
2
5.90066e-315 0
0
8 4-In OR~
219 675 315 0 5 22
0 14 23 24 18 11
0
0 0 1136 0
4 4072
-14 -24 14 -16
3 U8B
-3 -25 18 -17
1 b
-1 -45 6 -37
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 8 0
1 U
3311 0 0
2
5.90066e-315 0
0
14 Logic Display~
6 717 820 0 1 2
10 7
0
0 0 54368 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
7 check g
-25 -26 24 -18
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5736 0 0
2
44973.7 4
0
14 Logic Display~
6 719 741 0 1 2
10 8
0
0 0 54368 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
7 check f
-25 -26 24 -18
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3143 0 0
2
44973.7 5
0
14 Logic Display~
6 718 638 0 1 2
10 5
0
0 0 54368 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
7 check e
-25 -26 24 -18
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5835 0 0
2
44973.7 6
0
14 Logic Display~
6 738 505 0 1 2
10 9
0
0 0 54368 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
7 check d
-25 -26 24 -18
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5108 0 0
2
44973.7 7
0
14 Logic Display~
6 738 396 0 1 2
10 10
0
0 0 54368 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
7 check c
-25 -26 24 -18
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3320 0 0
2
44973.7 8
0
14 Logic Display~
6 738 296 0 1 2
10 11
0
0 0 54368 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
7 check b
-25 -26 24 -18
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
523 0 0
2
44973.7 9
0
8 4-In OR~
219 643 845 0 5 22
0 2 13 6 14 7
0
0 0 1136 0
4 4072
-14 -24 14 -16
3 U8A
-3 -25 18 -17
1 g
-2 -29 5 -21
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 8 0
1 U
3557 0 0
2
44973.7 10
0
5 4081~
219 509 810 0 3 22
0 16 15 19
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U5D
-12 -25 9 -17
3 B~D
-17 -25 4 -17
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
7246 0 0
2
44973.7 11
0
5 4081~
219 510 767 0 3 22
0 16 17 2
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U5C
-12 -25 9 -17
3 B~C
-12 -31 9 -23
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
3916 0 0
2
44973.7 12
0
5 4073~
219 510 615 0 4 22
0 16 17 3 20
0
0 0 1136 0
4 4073
-7 -24 21 -16
3 U6A
-12 -25 9 -17
4 B~CD
-17 -30 11 -22
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 6 0
1 U
614 0 0
2
44973.7 13
0
8 4-In OR~
219 617 543 0 5 22
0 14 13 4 6 21
0
0 0 1136 0
4 4072
-14 -24 14 -16
3 U2B
-3 -25 18 -17
7 4 terms
-23 -29 26 -21
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 2 0
1 U
8494 0 0
2
44973.7 14
0
5 4081~
219 510 550 0 3 22
0 22 15 6
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U5B
-12 -25 9 -17
3 C~D
-12 -31 9 -23
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
774 0 0
2
44973.7 15
0
5 4081~
219 508 491 0 3 22
0 23 22 13
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
3 ~BC
-12 -31 9 -23
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
715 0 0
2
44973.7 16
0
8 4-In OR~
219 675 180 0 5 22
0 14 22 4 25 12
0
0 0 1136 0
4 4072
-14 -24 14 -16
3 U2A
-3 -25 18 -17
1 a
-2 -29 5 -21
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
12 type:digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 2 0
1 U
3281 0 0
2
44973.7 17
0
5 4081~
219 510 326 0 3 22
0 22 3 24
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U3D
-12 -25 9 -17
2 CD
-9 -31 5 -23
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 3 0
1 U
3593 0 0
2
44973.7 18
0
5 4081~
219 511 383 0 3 22
0 17 15 18
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U3C
-12 -25 9 -17
4 ~C~D
-16 -31 12 -23
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
7233 0 0
2
44973.7 19
0
14 Logic Display~
6 740 161 0 1 2
10 12
0
0 0 54368 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
7 check a
-25 -26 24 -18
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3410 0 0
2
44973.7 20
0
5 4081~
219 510 228 0 3 22
0 16 3 25
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U3B
-12 -25 9 -17
2 BD
-11 -26 3 -18
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
3616 0 0
2
44973.7 21
0
5 4081~
219 510 168 0 3 22
0 23 15 4
0
0 0 1136 0
4 4081
-7 -24 21 -16
3 U3A
-12 -25 9 -17
4 ~B~D
-18 -31 10 -23
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
5202 0 0
2
44973.7 22
0
5 4049~
219 432 106 0 2 22
0 3 15
0
0 0 1136 270
4 4049
-7 -24 21 -16
3 U1C
16 -8 37 0
2 ~D
18 -9 32 -1
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 1 0
1 U
9145 0 0
2
44973.7 23
0
5 4049~
219 342 106 0 2 22
0 22 17
0
0 0 1136 270
4 4049
-7 -24 21 -16
3 U1B
16 -8 37 0
2 ~C
16 -7 30 1
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 1 0
1 U
9815 0 0
2
44973.7 24
0
5 4049~
219 255 105 0 2 22
0 16 23
0
0 0 1136 270
4 4049
-7 -24 21 -16
3 U1A
16 -8 37 0
2 ~B
15 -7 29 1
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
4766 0 0
2
44973.7 25
0
71
0 1 2 0 0 4096 0 0 17 29 0 3
558 752
558 832
626 832
2 0 3 0 0 4096 0 28 0 0 64 2
486 237
405 237
0 3 4 0 0 4112 0 0 21 56 0 3
573 185
573 548
600 548
3 1 5 0 0 12288 0 5 13 0 0 5
697 655
706 655
706 664
718 664
718 656
5 1 5 0 0 4224 0 6 13 0 0 4
993 153
993 657
718 657
718 656
2 0 6 0 0 8192 0 5 0 0 36 3
651 664
576 664
576 557
0 1 4 0 0 4224 0 0 5 56 0 3
557 185
557 646
651 646
7 0 7 0 0 4224 0 6 0 0 14 4
1005 153
1005 847
717 847
717 845
0 6 8 0 0 12416 0 0 6 15 0 4
719 756
719 757
999 757
999 153
0 4 9 0 0 12416 0 0 6 16 0 4
738 531
738 527
987 527
987 153
0 3 10 0 0 12416 0 0 6 17 0 4
737 422
737 418
981 418
981 153
0 2 11 0 0 8320 0 0 6 18 0 4
738 322
738 318
975 318
975 153
1 0 12 0 0 8320 0 6 0 0 19 4
969 153
969 184
740 184
740 187
5 1 7 0 0 0 0 17 11 0 0 3
676 845
717 845
717 838
5 1 8 0 0 0 0 7 12 0 0 3
698 756
719 756
719 759
3 1 9 0 0 0 0 8 14 0 0 5
708 522
726 522
726 531
738 531
738 523
5 1 10 0 0 0 0 9 15 0 0 5
708 414
726 414
726 422
738 422
738 414
5 1 11 0 0 0 0 10 16 0 0 5
708 315
726 315
726 322
738 322
738 314
5 1 12 0 0 0 0 24 27 0 0 5
708 180
728 180
728 187
740 187
740 179
0 2 13 0 0 4224 0 0 17 37 0 3
565 491
565 841
626 841
3 0 6 0 0 8320 0 17 0 0 36 3
626 850
550 850
550 550
4 0 14 0 0 4096 0 17 0 0 71 2
626 859
138 859
2 0 15 0 0 4096 0 18 0 0 63 2
485 819
435 819
1 0 16 0 0 4096 0 18 0 0 70 2
485 801
224 801
2 0 17 0 0 4096 0 19 0 0 65 2
486 776
345 776
1 0 16 0 0 4096 0 19 0 0 70 2
486 758
224 758
0 4 18 0 0 4224 0 0 7 47 0 3
582 329
582 770
648 770
3 3 19 0 0 4224 0 7 18 0 0 6
648 761
576 761
576 806
543 806
543 810
530 810
2 3 2 0 0 4224 0 7 19 0 0 4
648 752
539 752
539 767
531 767
1 0 14 0 0 8192 0 7 0 0 71 3
648 743
648 728
138 728
3 0 3 0 0 0 0 20 0 0 64 2
486 624
405 624
2 0 17 0 0 0 0 20 0 0 65 2
486 615
345 615
1 0 16 0 0 0 0 20 0 0 70 2
486 606
224 606
2 4 20 0 0 12416 0 8 20 0 0 4
662 531
653 531
653 615
531 615
1 5 21 0 0 8320 0 8 21 0 0 4
662 513
649 513
649 543
650 543
3 4 6 0 0 0 0 22 21 0 0 4
531 550
562 550
562 557
600 557
3 2 13 0 0 0 0 23 21 0 0 4
529 491
591 491
591 539
600 539
1 0 14 0 0 0 0 21 0 0 71 2
600 530
138 530
2 0 15 0 0 4096 0 22 0 0 63 2
486 559
435 559
1 0 22 0 0 4096 0 22 0 0 67 2
486 541
308 541
2 0 22 0 0 0 0 23 0 0 67 2
484 500
308 500
1 0 23 0 0 4096 0 23 0 0 68 4
484 482
263 482
263 483
258 483
4 0 3 0 0 4096 0 9 0 0 64 2
658 428
405 428
3 0 17 0 0 4096 0 9 0 0 65 2
658 419
345 419
2 0 16 0 0 4096 0 9 0 0 70 2
658 410
224 410
1 0 14 0 0 0 0 9 0 0 71 4
658 401
536 401
536 403
138 403
4 3 18 0 0 0 0 10 26 0 0 4
658 329
540 329
540 383
532 383
3 3 24 0 0 4224 0 10 25 0 0 4
658 320
539 320
539 326
531 326
2 0 15 0 0 4096 0 26 0 0 63 2
487 392
435 392
1 0 17 0 0 0 0 26 0 0 65 2
487 374
345 374
2 0 3 0 0 0 0 25 0 0 64 2
486 335
405 335
1 0 22 0 0 0 0 25 0 0 67 2
486 317
308 317
2 0 23 0 0 12288 0 10 0 0 68 4
658 311
541 311
541 280
258 280
1 0 14 0 0 0 0 10 0 0 71 4
658 302
550 302
550 259
138 259
4 3 25 0 0 4224 0 24 28 0 0 4
658 194
539 194
539 228
531 228
3 3 4 0 0 128 0 24 29 0 0 4
658 185
544 185
544 168
531 168
2 0 22 0 0 12288 0 24 0 0 67 4
658 176
551 176
551 147
308 147
1 0 14 0 0 0 0 24 0 0 71 4
658 167
558 167
558 135
138 135
1 0 16 0 0 0 0 28 0 0 70 2
486 219
224 219
1 0 23 0 0 0 0 29 0 0 68 2
486 159
258 159
2 0 15 0 0 0 0 29 0 0 63 2
486 177
435 177
1 0 3 0 0 0 0 30 0 0 64 2
435 88
405 88
2 0 15 0 0 4224 0 30 0 0 0 2
435 124
435 919
1 0 3 0 0 4224 0 1 0 0 0 2
405 80
405 920
2 0 17 0 0 4224 0 31 0 0 0 2
345 124
345 921
1 0 22 0 0 0 0 31 0 0 67 2
345 88
308 88
1 0 22 0 0 4224 0 3 0 0 0 2
308 80
308 923
2 0 23 0 0 4224 0 32 0 0 0 2
258 123
258 924
1 0 16 0 0 0 0 32 0 0 70 2
258 87
224 87
1 0 16 0 0 4224 0 2 0 0 0 2
224 81
224 926
1 0 14 0 0 4224 0 4 0 0 0 2
138 82
138 927
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
